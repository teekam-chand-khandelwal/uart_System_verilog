`include "uart_trans.sv"
`include "uart_gen.sv"
`include "uart_intf.sv"
`include "uart_driv.sv"
`include "uart_env.sv"
`include "uart_test.sv"
`include "tb_uart_top.sv"
